//拓展实验需要修改的代码部分很多，需要处理好每一个细节。指导教师提供的py程序、jpgtomif程序和字模生成软件给实验提供了很大帮助。
module lcd_display(
	input lcd_clk,
	input sys_rst_n,
	input[3:0]key,//对于按键控制问题，我们在输入端增加四个按键用于对屏幕展示内容的控制，并且注意，要在tcl文件中增加四行给四个按键分配引脚，分配与之前的实验相同
	input[10:0]pixel_xpos,
	input[10:0]pixel_ypos,
	output reg[15:0]pixel_data
	);
localparam PIC_X_START=11'd310;//原来的图片位置是屏幕左上角，这里修改为屏幕中心
localparam PIC_Y_START=11'd186;
localparam PIC_WIDTH=11'd180;//修改图片大小
localparam PIC_HEIGHT=11'd108;
localparam CHAR_X_START=11'd100;//原来的字也是放左上角，这里向中心移动了一点
localparam CHAR_Y_START=11'd100;
localparam CHAR_WIDTH=11'd256;//字符的宽、高，我们遇到了字符的宽不统一的问题（两个256一个352），最后将较短数组与96位0拼接，也就是在字符后加空格，统一了字符的宽
localparam CHAR_HEIGHT=11'd192;
localparam BACK_COLOR=16'hCE79;//修改背景颜色为浅灰色
localparam CHAR_COLOR=16'hF800;
localparam MODE_NAME=2'b00;//（四个模式：姓名、学号、学校、图片，对应0、1、2、3），处理按键输入转常驻模式信号的方式与流水灯拓展实验相同
localparam MODE_ID=2'b01;
localparam MODE_SCHOOL=2'b10;
localparam MODE_IMAGE=2'b11;
reg[14:0]rom_addr;//由于我们改变了图片的分辨率（从100*100的UCASLOGO改成180*108），这里的rom地址会出现越界问题，14位二进制不够用，最后生成的图片会发生上半部分重复出现下半部分不出现的问题，所以改成15位二进制解决问题
reg[3:0]key_last;//处理按键输入转常驻模式信号的方式与流水灯拓展实验相同
reg[1:0]mode;//处理按键输入转常驻模式信号的方式与流水灯拓展实验相同
reg[255:0]name_data[191:0];//我们使用了三个二维数组存储前三个字符屏幕画面，然后根据模式选择使用其中之一的数组
reg[255:0]id_data[95:0];
reg[351:0]school_data[31:0];
wire[351:0]current_char_line;//（这是选择的数组）
wire[10:0]char_x_pos;
wire[10:0]char_y_pos;
wire char_pixel;
wire rom_rd_en;
wire[15:0]rom_rd_data;
wire[3:0]key_pressed;//处理按键输入转常驻模式信号的方式与流水灯拓展实验相同
assign char_x_pos=pixel_xpos-CHAR_X_START;
assign char_y_pos=pixel_ypos-CHAR_Y_START;
assign rom_rd_en=1'b1;
assign key_pressed=(~key)&key_last;//处理按键输入转常驻模式信号的方式与流水灯拓展实验相同

always @(posedge lcd_clk or negedge sys_rst_n)begin//（对于这整个always逻辑），处理按键输入转常驻模式信号的方式与流水灯拓展实验相同
	if(!sys_rst_n)
		key_last<=4'b1111;
	else
		key_last<=key;
end
always @(posedge lcd_clk or negedge sys_rst_n)begin//（对于这整个always逻辑），按键信号转模式
	if(!sys_rst_n)
		mode<=MODE_NAME;
	else begin
		if(key_pressed[0])
			mode<=MODE_NAME;
		else if(key_pressed[1])
			mode<=MODE_ID;
		else if(key_pressed[2])
			mode<=MODE_SCHOOL;
		else if(key_pressed[3])
			mode<=MODE_IMAGE;
	end
end

assign current_char_line=(mode==MODE_NAME)?{96'b0,name_data[char_y_pos]}:(mode==MODE_ID)?{96'b0,id_data[char_y_pos]}:(mode==MODE_SCHOOL)?school_data[char_y_pos]:352'b0;//（同上）（这是选择的数组）
assign char_pixel=(char_x_pos<((mode==MODE_SCHOOL)?352:256))?current_char_line[((mode==MODE_SCHOOL)?352:256)-1-char_x_pos]:1'b0;

always @(posedge lcd_clk or negedge sys_rst_n)begin//（对于这整个always逻辑），关键修改：根据模式选择要输出的像素数据pixel_data
	if(!sys_rst_n)
		pixel_data<=BACK_COLOR;
	else if(mode==MODE_IMAGE)begin
		if((pixel_xpos>=PIC_X_START)&&(pixel_xpos<PIC_X_START+PIC_WIDTH)&&(pixel_ypos>=PIC_Y_START)&&(pixel_ypos<PIC_Y_START+PIC_HEIGHT))
			pixel_data<=rom_rd_data;
		else
			pixel_data<=BACK_COLOR;
	end
	else begin
		if((pixel_xpos>=CHAR_X_START)&&(pixel_xpos<CHAR_X_START+((mode==MODE_SCHOOL)?352:256))&&(pixel_ypos>=CHAR_Y_START)&&(pixel_ypos<CHAR_Y_START+((mode==MODE_NAME)?192:(mode==MODE_ID)?96:32)))
			pixel_data<=char_pixel?CHAR_COLOR:BACK_COLOR;
		else
			pixel_data<=BACK_COLOR;
	end
end
always @(posedge lcd_clk or negedge sys_rst_n)begin
	if(!sys_rst_n)
		rom_addr<=15'd0;
	else if((pixel_ypos>=PIC_Y_START)&&(pixel_ypos<PIC_Y_START+PIC_HEIGHT)&&(pixel_xpos>=PIC_X_START)&&(pixel_xpos<PIC_X_START+PIC_WIDTH))
		rom_addr<=rom_addr+1'b1;
	else if(pixel_ypos>=PIC_Y_START+PIC_HEIGHT)
		rom_addr<=15'd0;
end
rom_19440x16b u_rom_19440x16b(//注意，修改图片的过程，不仅要使用MegaWizard重新导入mif文件，还要在这里修改10000为19440，在这里遇到忘记修改的问题
	.address(rom_addr),
	.clock(lcd_clk),
	.rden(rom_rd_en),
	.q(rom_rd_data)
);
initial begin//（对于这整个initial逻辑），初始化这三个二维数组
	name_data[ 0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[ 1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[ 2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[ 3] <= 256'h0000000000000000000080000000000000000000000000000000000000000000;
	name_data[ 4] <= 256'h00000000000000000000E0000000000000000000000000000000000000000000;
	name_data[ 5] <= 256'h00000000000000000000F8000000000000000000000000000000000000000000;
	name_data[ 6] <= 256'h00000000000040000000F8000000008000000000000000000000000000000000;
	name_data[ 7] <= 256'h000000000000E0000000F000000001C000000000000000000000000000000000;
	name_data[ 8] <= 256'h007FFFFFFFFFF0000000F001FFFFFFE000000000000000000000000000000000;
	name_data[ 9] <= 256'h003FFFFFFFFFF8000000F000FFFFFFE000000000000000000000000000000000;
	name_data[10] <= 256'h0018003C0001E0000000F00061E003C000000000000000000000000000000000;
	name_data[11] <= 256'h0000003C0001E0000000F00001E0038000000000000000000000000000000000;
	name_data[12] <= 256'h0000003C0001E0000000F02001E0038000000000000000000000000000000000;
	name_data[13] <= 256'h0000003C0001E0000000F07001E0038000000000000000000000000000000000;
	name_data[14] <= 256'h0000003C0001E00007FFFFF801E0038000000000000000000000000000000000;
	name_data[15] <= 256'h0000003C0001E00003FFFFFC01E0038000000000000000000000000000000000;
	name_data[16] <= 256'h0000003C0001E0000100F00001E0038000000000000000000000000000000000;
	name_data[17] <= 256'h0000003C0001E0000000F00003C0078000000000000000000000000000000000;
	name_data[18] <= 256'h0000003C0001E1800000F00003C0078000000000000000000000000000000000;
	name_data[19] <= 256'h0000003C0001E3C00000F00003C0078000000000000000000000000000000000;
	name_data[20] <= 256'h0000003C0001E7E00000F0000780078000000000000000000000000000000000;
	name_data[21] <= 256'h0FFFFFFFFFFFFFF00000F0000780078000000000000000000000000000000000;
	name_data[22] <= 256'h07FFFFFFFFFFFFF80000F0000F00070000000000000000000000000000000000;
	name_data[23] <= 256'h030000380001E0000000F0000E060F0000000000000000000000000000000000;
	name_data[24] <= 256'h000000380001E0000000F0301E03FF0000000000000000000000000000000000;
	name_data[25] <= 256'h000000380001E0000000F0783C00FE0000000000000000000000000000000000;
	name_data[26] <= 256'h000000380001E0001FFFFFFC38003E0000000000000000000000000000000000;
	name_data[27] <= 256'h000000380001E0000FFFFFFE7000180000000000000000000000000000000000;
	name_data[28] <= 256'h000000780001E00004007001E000100000000000000000000000000000000000;
	name_data[29] <= 256'h000000780001E000000070038000000000000000000000000000000000000000;
	name_data[30] <= 256'h000000780001E000000070070000000000000000000000000000000000000000;
	name_data[31] <= 256'h000000780001E000000070042000020000000000000000000000000000000000;
	name_data[32] <= 256'h000000780001E000000070003800070000000000000000000000000000000000;
	name_data[33] <= 256'h000000780001E00000E070003FFFFF8000000000000000000000000000000000;
	name_data[34] <= 256'h007FFFFFFFFFE00000F870003FFFFFC000000000000000000000000000000000;
	name_data[35] <= 256'h003FFFFFFFFFE00000F870003C000F8000000000000000000000000000000000;
	name_data[36] <= 256'h001000700001E00000F070183C000F0000000000000000000000000000000000;
	name_data[37] <= 256'h000000F00001E00000F0703C3C000F0000000000000000000000000000000000;
	name_data[38] <= 256'h000000F00001E00000E07FFE3C000F0000000000000000000000000000000000;
	name_data[39] <= 256'h000000F00001000000E07FFF3C000F0000000000000000000000000000000000;
	name_data[40] <= 256'h000000E00000000000E070003C000F0000000000000000000000000000000000;
	name_data[41] <= 256'h000001E00000000000E070003C000F0000000000000000000000000000000000;
	name_data[42] <= 256'h000001E00000000000E070003C000F0000000000000000000000000000000000;
	name_data[43] <= 256'h000003C00000000000E070003C000F0000000000000000000000000000000000;
	name_data[44] <= 256'h000003C00000000001E070003C000F0000000000000000000000000000000000;
	name_data[45] <= 256'h000007800000000001E070003C000F0000000000000000000000000000000000;
	name_data[46] <= 256'h000007800000000001F070003C000F0000000000000000000000000000000000;
	name_data[47] <= 256'h00000F000000000001D870003FFFFF0000000000000000000000000000000000;
	name_data[48] <= 256'h00000E000000000001DC70003FFFFF0000000000000000000000000000000000;
	name_data[49] <= 256'h00001E000000000001CE70003C000F0000000000000000000000000000000000;
	name_data[50] <= 256'h00003C0000000000038770003C000F0000000000000000000000000000000000;
	name_data[51] <= 256'h00007800000000000383F0003C000E0000000000000000000000000000000000;
	name_data[52] <= 256'h0000F000000000000301F0003C00080000000000000000000000000000000000;
	name_data[53] <= 256'h0001E000000000000700F8003000000000000000000000000000000000000000;
	name_data[54] <= 256'h000380000000000006003F000000000000000000000000000000000000000000;
	name_data[55] <= 256'h000700000000000006001FF00000000000000000000000000000000000000000;
	name_data[56] <= 256'h001E0000000000000C0007FFF000000000000000000000000000000000000000;
	name_data[57] <= 256'h00380000000000000C0000FFFFFFFFF800000000000000000000000000000000;
	name_data[58] <= 256'h00E00000000000001800001FFFFFFFE000000000000000000000000000000000;
	name_data[59] <= 256'h0380000000000000100000007FFFFF8000000000000000000000000000000000;
	name_data[60] <= 256'h060000000000000020000000000FFF8000000000000000000000000000000000;
	name_data[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[64] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[65] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[66] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[67] <= 256'h0000000080000000000000000000000000000000000000000000000000000000;
	name_data[68] <= 256'h00000000E0000000000000C00000008000000000000000000000000000000000;
	name_data[69] <= 256'h00000000F8000000000001E0000003C000000000000000000000000000000000;
	name_data[70] <= 256'h00000400F80000001FFFFFF7FFFFFFE000000000000000000000000000000000;
	name_data[71] <= 256'h00000F00E00000000FFFFFFBFFFFFFF000000000000000000000000000000000;
	name_data[72] <= 256'h0FFFFF80E00000000603C0010078000000000000000000000000000000000000;
	name_data[73] <= 256'h07FFFF00E0001800000780000078000000000000000000000000000000000000;
	name_data[74] <= 256'h02000E00E0001C00000780000070000000000000000000000000000000000000;
	name_data[75] <= 256'h00000E00E0003E00000780000070000000000000000000000000000000000000;
	name_data[76] <= 256'h00000E00E0007E000007800000E0000000000000000000000000000000000000;
	name_data[77] <= 256'h00000E00E0007E000007000000E0000000000000000000000000000000000000;
	name_data[78] <= 256'h00000E00E000F800000F000000C0000000000000000000000000000000000000;
	name_data[79] <= 256'h00000E00E001F000000F000000C0000000000000000000000000000000000000;
	name_data[80] <= 256'h00000E00E003C000000E00000080020000000000000000000000000000000000;
	name_data[81] <= 256'h00000E00E0078000000E00018180070000000000000000000000000000000000;
	name_data[82] <= 256'h00000E00E00F0000001E0001FFFFFFC000000000000000000000000000000000;
	name_data[83] <= 256'h01000E00E01E0000001C0001FFFFFF8000000000000000000000000000000000;
	name_data[84] <= 256'h01800E00E03C0000001C0001E000070000000000000000000000000000000000;
	name_data[85] <= 256'h01FFFE00E0780000003C0001E000070000000000000000000000000000000000;
	name_data[86] <= 256'h01FFFE00E0E0000000380001E000070000000000000000000000000000000000;
	name_data[87] <= 256'h01E00E00E1C0000000380381E040070000000000000000000000000000000000;
	name_data[88] <= 256'h01E00F00E3800000007FFFC1E020070000000000000000000000000000000000;
	name_data[89] <= 256'h01C00800E6000000007FFFC1E038070000000000000000000000000000000000;
	name_data[90] <= 256'h01C00000EC00000000F80781E03E070000000000000000000000000000000000;
	name_data[91] <= 256'h01C00000F000010000F80781E03C070000000000000000000000000000000000;
	name_data[92] <= 256'h01C00000E000038000F80781E038070000000000000000000000000000000000;
	name_data[93] <= 256'h01C00000E00007C001F80781E078070000000000000000000000000000000000;
	name_data[94] <= 256'h01C003FFFFFFFFE001B80781E078070000000000000000000000000000000000;
	name_data[95] <= 256'h03C011FFFFFFFFF003B80781E078070000000000000000000000000000000000;
	name_data[96] <= 256'h03C01CC0E080000003380781E078070000000000000000000000000000000000;
	name_data[97] <= 256'h07FFFE00E080000006380781E078070000000000000000000000000000000000;
	name_data[98] <= 256'h07FFFE00E0C0000004380781E078070000000000000000000000000000000000;
	name_data[99] <= 256'h03803C00E0C000000C380781E078070000000000000000000000000000000000;
	name_data[100] <= 256'h01003800E060000018380781E078070000000000000000000000000000000000;
	name_data[101] <= 256'h00003800E060000010380781E078070000000000000000000000000000000000;
	name_data[102] <= 256'h00003800E070000000380781E070070000000000000000000000000000000000;
	name_data[103] <= 256'h00003800E030000000380781E070070000000000000000000000000000000000;
	name_data[104] <= 256'h00003800E038000000380781E0F0070000000000000000000000000000000000;
	name_data[105] <= 256'h00003800E038000000380781E0F0070000000000000000000000000000000000;
	name_data[106] <= 256'h00003800E01C000000380781E0F0070000000000000000000000000000000000;
	name_data[107] <= 256'h00003800E01E000000380781E0E0070000000000000000000000000000000000;
	name_data[108] <= 256'h00003800E00E0000003FFF81E1E0060000000000000000000000000000000000;
	name_data[109] <= 256'h00007800E0070000003FFF8181E0040000000000000000000000000000000000;
	name_data[110] <= 256'h00007800E00780000038078003C6000000000000000000000000000000000000;
	name_data[111] <= 256'h00007800E003C0000038078003C3800000000000000000000000000000000000;
	name_data[112] <= 256'h00007000E003E000003807000781E00000000000000000000000000000000000;
	name_data[113] <= 256'h00007000E001F000003804000F00F80000000000000000000000000000000000;
	name_data[114] <= 256'h00007000E018F800003800000F003E0000000000000000000000000000000000;
	name_data[115] <= 256'h0000F000E0607E00003800001E001F0000000000000000000000000000000000;
	name_data[116] <= 256'h0000F000E1C03F80003800007C000FC000000000000000000000000000000000;
	name_data[117] <= 256'h0000E000E7803FE000200000F8000FC000000000000000000000000000000000;
	name_data[118] <= 256'h03C1E000FF001FF800000001E00007E000000000000000000000000000000000;
	name_data[119] <= 256'h00FFE000FE000FE000000007C00003E000000000000000000000000000000000;
	name_data[120] <= 256'h003FC001FC0007800000000F000001E000000000000000000000000000000000;
	name_data[121] <= 256'h001F8001F80001000000003C000001E000000000000000000000000000000000;
	name_data[122] <= 256'h001F0000F0000000000000F0000000E000000000000000000000000000000000;
	name_data[123] <= 256'h000E000060000000000003800000004000000000000000000000000000000000;
	name_data[124] <= 256'h000000000000000000000C000000000000000000000000000000000000000000;
	name_data[125] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[126] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[127] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[128] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[129] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[130] <= 256'h0000000200000000000000000000000000080000000000000000000000000000;
	name_data[131] <= 256'h00000003800000000000000000000000000E0000000000000000000000000000;
	name_data[132] <= 256'h00000003E00000000000000000000000000F8000000000000000000000000000;
	name_data[133] <= 256'h00000003E00000000000000000000200000F8000000000000000000000000000;
	name_data[134] <= 256'h00000003C00000000000000000000700000F0000000002000000000000000000;
	name_data[135] <= 256'h00000003800000000000000000000F80000E0000000007000000000000000000;
	name_data[136] <= 256'h000000038000020007FFFFFFFFFFFFC0000E000000000F800000000000000000;
	name_data[137] <= 256'h000000038000070003FFFFFFFFFFFFE0000E01FFFFFFFFC00000000000000000;
	name_data[138] <= 256'h0000000380000F800100000380000000000E00FFFFFFFFE00000000000000000;
	name_data[139] <= 256'h0FFFFFFFFFFFFFC00000000380000000000E0040000000000000000000000000;
	name_data[140] <= 256'h07FFFFFFFFFFFFE00000000380000000000E0000000000000000000000000000;
	name_data[141] <= 256'h0300007B900000000000000380000000000E0000000000000000000000000000;
	name_data[142] <= 256'h0000007B980000000000000380000000000F0000000000000000000000000000;
	name_data[143] <= 256'h000000F38C0000000000000380000000000FC000000000000000000000000000;
	name_data[144] <= 256'h000001E38E0000000000000380000000000EF000000000000000000000000000;
	name_data[145] <= 256'h000003C3860000000040000380001000000E7810000020000000000000000000;
	name_data[146] <= 256'h00000383830000000020000380003C00010E3C18000070000000000000000000;
	name_data[147] <= 256'h0000078383800000003FFFFFFFFFFE00010E3E1FFFFFFC000000000000000000;
	name_data[148] <= 256'h00000F0381E00000003FFFFFFFFFFE00010E1E1FFFFFFE000000000000000000;
	name_data[149] <= 256'h00001E0380F000000038000380003C00010E1E1E000078000000000000000000;
	name_data[150] <= 256'h00003803807C00000038000380003C00030E0E1E000078000000000000000000;
	name_data[151] <= 256'h00007003803E00000038000380003C00030E0E1E000078000000000000000000;
	name_data[152] <= 256'h0000E003801FC0000038000380003C00030E041E000078000000000000000000;
	name_data[153] <= 256'h0001C003800FF000003870038E003C00070E001E000078000000000000000000;
	name_data[154] <= 256'h000780038007FE0000383C0387803C00070E001E000078000000000000000000;
	name_data[155] <= 256'h000E00020021FFF000381E0383E03C000F0E001E000078000000000000000000;
	name_data[156] <= 256'h001C00000070FFF000380F8381F03C001F0E001E000078000000000000000000;
	name_data[157] <= 256'h0070FFFFFFF83F8000380F8380F83C003F0E001E000078000000000000000000;
	name_data[158] <= 256'h00C07FFFFFFC0E00003807C380783C003E0E001FFFFFF8000000000000000000;
	name_data[159] <= 256'h0380000000FE0200003803C380383C00000E001FFFFFF8000000000000000000;
	name_data[160] <= 256'h0E00000001F800000038038380383C00000E001E000078000000000000000000;
	name_data[161] <= 256'h1800000003C000000038018380183C00000E001E000078000000000000000000;
	name_data[162] <= 256'h00000000070000000038000380003C00000E001E000078000000000000000000;
	name_data[163] <= 256'h000000011C0000000038000380003C00000E001E000078000000000000000000;
	name_data[164] <= 256'h00000001F80000000038000380003C00000E001E000078000000000000000000;
	name_data[165] <= 256'h00000001E00000000038000380003C00000E001E000078000000000000000000;
	name_data[166] <= 256'h00000001F80000000038000380003C00000E001E000078000000000000000000;
	name_data[167] <= 256'h00000001F00001000038E00380003C00000E001E000078000000000000000000;
	name_data[168] <= 256'h00000001E00003800038780386003C00000E001E000078000000000000000000;
	name_data[169] <= 256'h00000001E00007C000383E0383C03C00000E001E000078000000000000000000;
	name_data[170] <= 256'h0FFFFFFFFFFFFFE000381F0381F03C00000E001E000078000000000000000000;
	name_data[171] <= 256'h07FFFFFFFFFFFFF000380F8380F83C00000E001FFFFFF8000000000000000000;
	name_data[172] <= 256'h02000001E00000000038078380783C00000E001FFFFFF8000000000000000000;
	name_data[173] <= 256'h00000001E000000000380783807C3C00000E001E000078000000000000000000;
	name_data[174] <= 256'h00000001E000000000380383803C3C00000E001E000078000000000000000000;
	name_data[175] <= 256'h00000001E00000000038030380183C00000E001E000070000000000000000000;
	name_data[176] <= 256'h00000001E00000000038000380183C00000E001C000040000000000000000000;
	name_data[177] <= 256'h00000001E00000000038000380003C00000E0010000000000000000000000000;
	name_data[178] <= 256'h00000001E00000000038000380003C00000E0000000000000000000000000000;
	name_data[179] <= 256'h00000001E00000000038000380003C00000E0000000001800000000000000000;
	name_data[180] <= 256'h00000001E00000000038000380003C00000E0000000003C00000000000000000;
	name_data[181] <= 256'h00000001E00000000038000380007800000E0000000007E00000000000000000;
	name_data[182] <= 256'h00000601E00000000038000380FFF800000E1FFFFFFFFFF00000000000000000;
	name_data[183] <= 256'h000007FFE000000000380003800FF800000E0FFFFFFFFFF80000000000000000;
	name_data[184] <= 256'h0000007FC0000000003800038003F800000E0400000000000000000000000000;
	name_data[185] <= 256'h0000001FC0000000003800030001F000000E0000000000000000000000000000;
	name_data[186] <= 256'h0000000F80000000003000040000E000000E0000000000000000000000000000;
	name_data[187] <= 256'h00000007000000000040000000008000000F0000000000000000000000000000;
	name_data[188] <= 256'h0000000400000000000000000000000000080000000000000000000000000000;
	name_data[189] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[190] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	name_data[191] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 3] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 4] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 5] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[ 6] <= 256'h07E003C007E007C07E7C07E003C003C007C007C007E001E003C003C007C00000;
	id_data[ 7] <= 256'h083806200838186018300C300620062018201820083806180620062018600000;
	id_data[ 8] <= 256'h10180C3010183030182018180C300C303010301010180C180C300C3030300000;
	id_data[ 9] <= 256'h200C1818200C30181860300C1818181830183018200C08181818181830180000;
	id_data[10] <= 256'h200C1818200C30181840300C1818181860086008200C18001818181830180000;
	id_data[11] <= 256'h300C1808300C30181880300C18081808600C600C300C10001808180830180000;
	id_data[12] <= 256'h300C300C300C00181880380C300C300C600C600C300C1000300C300C00180000;
	id_data[13] <= 256'h000C300C000C001819003808300C300C600C600C000C3000300C300C00180000;
	id_data[14] <= 256'h0018300C0018003019001E18300C300C600C600C001833E0300C300C00300000;
	id_data[15] <= 256'h0018300C001800601B000F20300C300C600C600C00183630300C300C00600000;
	id_data[16] <= 256'h0030300C003003C01D8007C0300C300C701C701C00303818300C300C03C00000;
	id_data[17] <= 256'h0060300C006000701D8018F0300C300C302C302C00603808300C300C00700000;
	id_data[18] <= 256'h00C0300C00C0001818C03078300C300C186C186C00C0300C300C300C00180000;
	id_data[19] <= 256'h0180300C0180000818C03038300C300C0F8C0F8C0180300C300C300C00080000;
	id_data[20] <= 256'h0300300C0300000C1860601C300C300C000C000C0300300C300C300C000C0000;
	id_data[21] <= 256'h0200300C0200000C1860600C300C300C001800180200300C300C300C000C0000;
	id_data[22] <= 256'h040418080404300C1830600C18081808001800180404300C18081808300C0000;
	id_data[23] <= 256'h080418180804300C1830600C18181818001000100804180C18181818300C0000;
	id_data[24] <= 256'h10041818100430081830600C1818181830303030100418081818181830080000;
	id_data[25] <= 256'h200C0C30200C3018181830180C300C3030603060200C0C180C300C3030180000;
	id_data[26] <= 256'h3FF806203FF81830181818300620062030C030C03FF80E300620062018300000;
	id_data[27] <= 256'h3FF803C03FF807C07E3E07C003C003C00F800F803FF803E003C003C007C00000;
	id_data[28] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[29] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[30] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[31] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[32] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[33] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[34] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[35] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[36] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[37] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[38] <= 256'h0FF003C007E007C07E7C07E003C003C007C007C007E001E003C007E007C00000;
	id_data[39] <= 256'h1E7806200838186018300C300620062018201820083806180620083818200000;
	id_data[40] <= 256'h383C0C3010183030182018180C300C303010301010180C180C30101830100000;
	id_data[41] <= 256'h381C1818200C30181860300C1818181830183018200C08181818200C30180000;
	id_data[42] <= 256'h781C1818200C30181840300C1818181860086008200C18001818200C60080000;
	id_data[43] <= 256'h781C1808300C30181880300C18081808600C600C300C10001808300C600C0000;
	id_data[44] <= 256'h7C1C300C300C00181880380C300C300C600C600C300C1000300C300C600C0000;
	id_data[45] <= 256'h381C300C000C001819003808300C300C600C600C000C3000300C000C600C0000;
	id_data[46] <= 256'h003C300C0018003019001E18300C300C600C600C001833E0300C0018600C0000;
	id_data[47] <= 256'h0038300C001800601B000F20300C300C600C600C00183630300C0018600C0000;
	id_data[48] <= 256'h0070300C003003C01D8007C0300C300C701C701C00303818300C0030701C0000;
	id_data[49] <= 256'h00F0300C006000701D8018F0300C300C302C302C00603808300C0060302C0000;
	id_data[50] <= 256'h01E0300C00C0001818C03078300C300C186C186C00C0300C300C00C0186C0000;
	id_data[51] <= 256'h03C0300C0180000818C03038300C300C0F8C0F8C0180300C300C01800F8C0000;
	id_data[52] <= 256'h0780300C0300000C1860601C300C300C000C000C0300300C300C0300000C0000;
	id_data[53] <= 256'h0F00300C0200000C1860600C300C300C001800180200300C300C020000180000;
	id_data[54] <= 256'h0E0618080404300C1830600C18081808001800180404300C1808040400180000;
	id_data[55] <= 256'h1C0E18180804300C1830600C18181818001000100804180C1818080400100000;
	id_data[56] <= 256'h380C1818100430081830600C1818181830303030100418081818100430300000;
	id_data[57] <= 256'h701C0C30200C3018181830180C300C3030603060200C0C180C30200C30600000;
	id_data[58] <= 256'h7FFC06203FF81830181818300620062030C030C03FF80E3006203FF830C00000;
	id_data[59] <= 256'h7FFC03C03FF807C07E3E07C003C003C00F800F803FF803E003C03FF80F800000;
	id_data[60] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[61] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[64] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[65] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[66] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[67] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[68] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[69] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[70] <= 256'h0FF003C007E007C07E7C07E003C003C007C007C003C001E003C007E003C00000;
	id_data[71] <= 256'h1E7806200838186018300C300620062018201820062006180620083806200000;
	id_data[72] <= 256'h383C0C3010183030182018180C300C30301030100C300C180C3010180C300000;
	id_data[73] <= 256'h381C1818200C30181860300C1818181830183018181808181818200C18180000;
	id_data[74] <= 256'h781C1818200C30181840300C1818181860086008181818001818200C18180000;
	id_data[75] <= 256'h781C1808300C30181880300C18081808600C600C180810001808300C18080000;
	id_data[76] <= 256'h7C1C300C300C00181880380C300C300C600C600C300C1000300C300C300C0000;
	id_data[77] <= 256'h381C300C000C001819003808300C300C600C600C300C3000300C000C300C0000;
	id_data[78] <= 256'h003C300C0018003019001E18300C300C600C600C300C33E0300C0018300C0000;
	id_data[79] <= 256'h0038300C001800601B000F20300C300C600C600C300C3630300C0018300C0000;
	id_data[80] <= 256'h0070300C003003C01D8007C0300C300C701C701C300C3818300C0030300C0000;
	id_data[81] <= 256'h00F0300C006000701D8018F0300C300C302C302C300C3808300C0060300C0000;
	id_data[82] <= 256'h01E0300C00C0001818C03078300C300C186C186C300C300C300C00C0300C0000;
	id_data[83] <= 256'h03C0300C0180000818C03038300C300C0F8C0F8C300C300C300C0180300C0000;
	id_data[84] <= 256'h0780300C0300000C1860601C300C300C000C000C300C300C300C0300300C0000;
	id_data[85] <= 256'h0F00300C0200000C1860600C300C300C00180018300C300C300C0200300C0000;
	id_data[86] <= 256'h0E0618080404300C1830600C18081808001800181808300C1808040418080000;
	id_data[87] <= 256'h1C0E18180804300C1830600C18181818001000101818180C1818080418180000;
	id_data[88] <= 256'h380C1818100430081830600C1818181830303030181818081818100418180000;
	id_data[89] <= 256'h701C0C30200C3018181830180C300C30306030600C300C180C30200C0C300000;
	id_data[90] <= 256'h7FFC06203FF81830181818300620062030C030C006200E3006203FF806200000;
	id_data[91] <= 256'h7FFC03C03FF807C07E3E07C003C003C00F800F8003C003E003C03FF803C00000;
	id_data[92] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[93] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[94] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	id_data[95] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
	school_data[ 0] <= 352'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	school_data[ 1] <= 352'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	school_data[ 2] <= 352'h0003800008000020000000800004010000002000000100000004010000600800000600000002000000002000;
	school_data[ 3] <= 352'h0003C0000FFFFFF8000C00E00102018010201800000180000102018000700E00000300000003800000003800;
	school_data[ 4] <= 352'h000380000C000030003C00C0018303801FF00C0000018000018303800C618C00000180000003000000103000;
	school_data[ 5] <= 352'h000380000C00003007E000C000C38300186408100001800000C38300066318000001C000000300000FFC6020;
	school_data[ 6] <= 352'h000380000C00033038C000C000E186001867FFF80001800000E1860007661800040080100003000008187FF0;
	school_data[ 7] <= 352'h000380000CFFFFB000C060C0006184001844003000018000006184000264100007FFFFF80403008008184060;
	school_data[ 8] <= 352'h0C0380700C01803000C030C000610C0018CC00200001801000610C00006910080400003007FFFFC00818C0C0;
	school_data[ 9] <= 352'h0FFFFFF80C01803000C018C000400818188C004000018038004008183FFFFFFC0C000060060300C00818A0C0;
	school_data[10] <= 352'h0E0380700C01803000C018C00FFFFFFC188000003FFFFFFC0FFFFFFC00E030600C000040060300C008199180;
	school_data[11] <= 352'h0E0380700C01803000C400C00C00001819000180000180000C00001801F8306018000200060300C008191100;
	school_data[12] <= 352'h0E0380700C0180303FFE00C00C0000301903FFC0000180000C000030016E706001FFFF00060300C00FFA0B00;
	school_data[13] <= 352'h0E0380700C01843000C000C01C00024018800000000380001C0002400266506000000700060300C009920E00;
	school_data[14] <= 352'h0E0380700C7FFE3000C040C019FFFF00184000000003800019FFFF000462904000001C0007FFFFC001800F00;
	school_data[15] <= 352'h0E0380700C01803001C060C0000007001860003000034000000007001860904000003000060300C001801B80;
	school_data[16] <= 352'h0E0380700C01A03001F030C000001C00182FFFF00003400000001C00204108C000014000060300C0119030E0;
	school_data[17] <= 352'h0E0380700C01983003DC10C00000300018304600000320000000300000E008C000018000060300C01DF8607C;
	school_data[18] <= 352'h0FFFFFF00C018C3002CC00CC0001400018304600000620000001400000C208C000018018060300C01980C058;
	school_data[19] <= 352'h0E0380700C018E3006C400FC000180101830460000063000000180103FFF0C803FFFFFFC060300C019837FF8;
	school_data[20] <= 352'h0E0380700C01843004C40FC00001803818304600000610000001803801860D8000018000060300C0198C4060;
	school_data[21] <= 352'h080380000C01843008C1F0C03FFFFFFC19E0C600000C08003FFFFFFC010605800001800007FFFFC019804060;
	school_data[22] <= 352'h000380000C01833010C600C00001800018C0C600000C0C0000018000030C070000018000060300C019804060;
	school_data[23] <= 352'h000380000DFFFFB020C000C000018000180086080018060000018000038C0700000180000603000819804060;
	school_data[24] <= 352'h000380000C00003040C000C00001800018018608003003000001800000780700000180000003000819B84060;
	school_data[25] <= 352'h000380000C00003000C000C000018000180186080060038000018000003F0D8000018000000300081BC04060;
	school_data[26] <= 352'h000380000C00003000C000C0000180001803060800C001E00001800000E318E000018000000300083E004060;
	school_data[27] <= 352'h000380000FFFFFF000C000C00001800018060608018000F80001800001813070000180000003001838007FE0;
	school_data[28] <= 352'h000380000C00003000C000C0001F80001808071C06000038001F80000600C03E003F80000003FFFC00004060;
	school_data[29] <= 352'h000380000C00003000C000C000078000187003F8180000100007800038010010000780000001FFF800004060;
	school_data[30] <= 352'h0003800008000000008000800002000010000000200000000002000000060000000200000000000000000000;
	school_data[31] <= 352'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end
endmodule